`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Portland State University, ECE 540 Embedded System
// Project 2: RoJobot world
// Copyright by Dung Le
//
// Module Name:    Icon 
// Create Date:    15:00:42 10/31/2012 
// Target Devices: nexys 3 
// Tool versions: ISE 14.2
//
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments:  
//
//////////////////////////////////////////////////////////////////////////////////
module Icon(
	//
	////////////////////////////////////////////////////////////////////////////
	// INPUT
	////////////////////////////////////////////////////////////////////////////
	//
	input        clk, 
	input [7:0]  LocX,	
	input [7:0]  LocY,
	input [7:0]  BotInfo,
	input [9:0]  pixel_row, pixel_col,
	//
	////////////////////////////////////////////////////////////////////////////
	// OUTPUT
	////////////////////////////////////////////////////////////////////////////
	//
	output reg [7:0] icon
	);
	//
	////////////////////////////////////////////////////////////////////////////
	// SIGNALS
	////////////////////////////////////////////////////////////////////////////	
	//
	// remapping robot location to VGA display resolution
	wire [9:0] robot_disp_locX, robot_disp_locY;	
	// position of image's left top conner pixel
	reg [9:0] robot_icon_start_pixel_X;
	reg [9:0] robot_icon_start_pixel_Y;
	reg [8:0] pixel_address; // currently design to have 2 images (256 byte each) in ROM
	reg enable;
	wire [7:0] pixel_out;    // pixel getting from rom
	// x and y indexing into rom image
	reg [3:0] x,y;
	//
	////////////////////////////////////////////////////////////////////////////
	// Instantiate robot Icon ROM (generated by Xilinx Core Gnerator)
	////////////////////////////////////////////////////////////////////////////
	//
	icon_rom rb(
	.clka(clk),
	//.ena(enable),
	.addra(pixel_address),
	.douta(pixel_out)
	);
	//
	////////////////////////////////////////////////////////////////////////////
	// Start of module logic 
	////////////////////////////////////////////////////////////////////////////
	//
	// mapping 128x128 world to 512x512 display image
	//
	assign robot_disp_locX = {LocX,2'b00};
	assign robot_disp_locY = {LocY,2'b00};
	//
	// calculate icon start pixel position (left conner)
	//	
	always @( posedge clk) begin
		if (LocX == 8'b0 || LocX == 8'b1)
			robot_icon_start_pixel_X <= 10'b0;			           // clipping if robot at boundary
		else
			robot_icon_start_pixel_X <= robot_disp_locX - 10'd6; // line center alignment
	end
	//
	always @( posedge clk) begin
		if (LocY == 8'b0 || LocY == 8'b1)
			robot_icon_start_pixel_Y <= 10'b0;			
		else
			robot_icon_start_pixel_Y <= robot_disp_locY - 10'd6; 
	end
	//
	// calculate rom indexes using current pixel[row][col] and icon's left top conner pixel
	//
	always @ (posedge clk) begin
		y <= pixel_row[3:0] - robot_icon_start_pixel_Y[3:0];
		x <= pixel_col[3:0] - robot_icon_start_pixel_X[3:0];
	end
	//
	// Pixel Address transformation,
	// whenever row and col addr fall into the 16x16 area occupied by robot icon
	//	
	always @ (posedge clk) begin
		if( pixel_col >= robot_icon_start_pixel_X  
		&& pixel_col <= (robot_icon_start_pixel_X + 10'd15)
		&& pixel_row >= robot_icon_start_pixel_Y
		&& pixel_row <= (robot_icon_start_pixel_Y + 10'd15)
		) 
		begin
			//
		   // Indexing icon in ROM:
			// + first image: lower 256 bytes, orientation is 0 degree (North)
			// + second image: upper 256 bytes, orientation is 45 degree (North East)
			//
			// Image transformation: 
			// image[y][x]                   /* assuming this is the original orientation */
			// image[original_height - x][y] /* 90 degrees cw */
			// image[x][original_width - y]  /* rotated 90 degrees ccw */
			// image[original_height - y][original_width - x] /* 180 degrees */
			//
			case (BotInfo[2:0])
				// 0 degree. use first image
				3'd0:	pixel_address <= {1'b0, y, x};
				
				// 45 degree, use second image
				3'd1:	pixel_address <= {1'b1, y, x};
				
				// 90 degree, use first image, indexing rom[height - x][y]
				3'd2:	pixel_address <= {1'b0, 4'b1111 - x, y};
				
				// 135 degree, use second image, indexing rom[height - x][y]
				3'd3:	pixel_address <= {1'b1, 4'b1111 - x, y};
				
				// 180 degree, use first image, indexing rom[height - y][width - x]
				3'd4:	pixel_address <= {1'b0,4'b1111 - y, 4'b1111 - x};
				
				// 225 degree, use second image, indexing rom[height - y][width - x]
				3'd5:	pixel_address <= {1'b1,4'b1111 - y, 4'b1111 - x};
				
				// 270 degree, use first image, indexing rom[x][width - y]
				3'd6:	pixel_address <= {1'b0, x, 4'b1111 - y};	
				
				// 315 degree, use second image, indexing rom[x][width - y]
				3'd7:	pixel_address <= {1'b1, x, 4'b1111 - y};			
			endcase
			// get RGB byte from icon_rom
			icon <= pixel_out;  
		end
		else begin
			pixel_address <= 0;
			icon <= 0;	        // 0 means transparent
		end
	end
	
endmodule

